*$
**************** Power Discrete MOSFET Electrical Circuit Model *****************
** Product Name: FDPF3N50NZ 
** 500V N-Channel MOSFET and TO-220F
** Model Type: BSIM3V3
**-------------------------------------------------------------------------------
.SUBCKT FDPF3N50NZ 2 1 3    
*Nom Temp=25 deg C
Dbody 7 5    DbodyMOD
Dbreak 5 11  DbreakMOD
Ebreak 11 7 17 7 500
Lgate 1 9    1.474e-9
Ldrain 2 5   1.474e-9
Lsource 3 7  9.664e-10
RLgate 1 9   14.74
RLdrain 2 5  14.74
RLsource 3 7 9.664
Rgate 9 6    0.5
It 7 17      1
Rbreak 17 7  RbreakMOD 1
.MODEL RbreakMOD RES (TC1=1.08e-3 TC2=-1.12e-6)
.MODEL DbodyMOD D (IS=1.45e-13  N=1.0     RS=2.64e-2   TRS1=2.75e-3   TRS2=1.5e-6 
+ CJO=2.76e-10     M=0.62       VJ=0.72   TT=2.16e-7   XTI=3          EG=1.18)
.MODEL DbreakMOD D (RS=100e-3 TRS1=1.0e-3 TRS2=5.0e-6)
Rdrain 5 16 RdrainMOD 2.1
.MODEL RdrainMOD RES (TC1=8.45e-3 TC2=2.16e-5)
D_ZENER 7 9 Dzener
.MODEL Dzener D (IS=1e-12 N=2.0 BV=45.0 IBV=2.5e-4)
M_BSIM3 16 6 7 7 Bsim3 W=0.504 L=2.0e-6 NRS=1
.MODEL Bsim3 NMOS (LEVEL=7 VERSION=3.1 MOBMOD=3 CAPMOD=2 PARAMCHK=1 NQSMOD=0
+ TOX=1100e-10    XJ=1.4e-6      NCH=1.43e17
+ U0=700          VSAT=2.5e5     DROUT=1.0
+ DELTA=0.1       PSCBE2=0       RSH=1.19e-3
+ VTH0=4.18       VOFF=-0.1      NFACTOR=1.1
+ LINT=3.0e-7     DLC=3.0e-7     FC=0.5
+ CGSO=1.05e-15   CGSL=0         CGDO=2.25e-12  
+ CGDL=3.85e-10   CJ=0           CF=0
+ CKAPPA=0.2      KT1=-2.27      KT2=0
+ UA1=3.0e-9      NJ=10)
.ENDS
*$
******************** Power Discrete MOSFET Thermal Model ************************
** 500V N-Channel MOSFET and TO-220F
**-------------------------------------------------------------------------------
.SUBCKT FDPF3N50NZ_Thermal TH TL
CTHERM1 TH 6 2.04e-5
CTHERM2 6 5  1.14e-3
CTHERM3 5 4  2.82e-3
CTHERM4 4 3  3.64e-3
CTHERM5 3 2  8.02e-3
CTHERM6 2 TL 3.12e-2
RTHERM1 TH 6 2.00e-2
RTHERM2 6 5  1.20e-1
RTHERM3 5 4  2.60e-1
RTHERM4 4 3  3.60e-1
RTHERM5 3 2  8.10e-1
RTHERM6 2 TL 3.03e+0
.ENDS FDPF3N50NZ_Thermal
**-------------------------------------------------------------------------------
** Creation: Oct.-21-2015   Rev.: 0.0
** Fairchild Semiconductor
*$

