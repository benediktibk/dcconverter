**************** Power Discrete MOSFET Electrical Circuit Model *****************
** Product Name: FQP3P50
** 500V P-Channel MOSFET
** Model Type: BSIM3V3
**-------------------------------------------------------------------------------
.SUBCKT FQP3P50 2 1 3    
*Nom Temp=25 deg C
Dbody 5 7 DbodyMOD
Dbreak 7 11 DbreakMOD
Lgate 1 9 1.125e-9
Ldrain 2 5 5.00e-10
Lsource 3 7 9.66e-10
RLgate 1 9 11.25
RLdrain 2 5 5.00
RLsource 3 7 9.66
Rgate 9 6 0.5
It 7 17 1
Ebreak 5 11 17 7 -500
Rbreak 17 7 RbreakMOD 1
.MODEL RbreakMOD RES (TC1=8.2e-4 TC2=-1.05e-6)
.MODEL DbodyMOD D (IS=1.08e-15  N=1.0    RS=0.152   TRS1=1.0e-6  TRS2=1.1e-7
+ CJO=6.52e-10     M=0.42       VJ=0.65  TT=4.39e-7 XTI=3        EG=1.24)
.MODEL DbreakMOD D (RS=0.1 TRS1=1e-3 TRS2=1e-6)
Rdrain 5 16 RdrainMOD 3.9
.MODEL RdrainMOD RES (TC1=7.31e-3 TC2=1.14e-5)
M_BSIM3 16 6 7 7 Bsim3 W=0.86 L=2.0e-6 NRS=1
.MODEL Bsim3 PMOS (LEVEL=7 VERSION=3.1 MOBMOD=3 CAPMOD=2 PARAMCHK=1 NQSMOD=0
+ TOX=970e-10      XJ=1.0e-6       NCH=1.1e17
+ U0=250           VSAT=5.0e5      DROUT=1.0
+ DELTA=0.1        PSCBE2=0        RSH=1.5e-3
+ VTH0=-3.55       VOFF=-0.1       NFACTOR=1.1     
+ LINT=2.7e-8      DLC=2.7e-8      CGSO=1.1e-15
+ CGSL=0           CGDO=6.5e-15    CGDL=7.82e-10
+ CJ=0             CF=0            CKAPPA=0.2
+ KT1=-1.08        KT2=0           UA1=-7.2e-9
+ NJ=10            FC=0.5)
.ENDS

******************* Power Discrete MOSFET Thermal Model ************************
** Product: FQP3P50
** Package: TO-220
**------------------------------------------------------------------------------
.SUBCKT FQP3P50_THERMAL TH TL
CTHERM1 TH 6 8.04e-4
CTHERM2 6 5  4.28e-3
CTHERM3 5 4  8.34e-3
CTHERM4 4 3  1.62e-2
CTHERM5 3 2  2.02e-1
CTHERM6 2 TL 5.42e-1
RTHERM1 TH 6 1.30e-2
RTHERM2 6 5  2.88e-2
RTHERM3 5 4  3.68e-2
RTHERM4 4 3  4.12e-1
RTHERM5 3 2  4.41e-1
RTHERM6 2 TL 5.38e-1
.ENDS FQP3P50_THERMAL
**-----------------------------------------------------------------------------
** Creation: Mar.-16-2012   Rev.:0.0
** Fairchild Semiconductor

