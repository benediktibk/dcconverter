*$
****************** Power Discrete MOSFET Electrical Circuit Model *******************
** Product Name: FQB1P50
** 500V P-Channel MOSFET
** Model Type: BSIM3V3
**----------------------------------------------------------------------------------
.subckt FQB1P50 2 1 3
*Nom Temp=25 deg C
Dbody 5 7 DbodyMOD
Dbreak 7 11 DbreakMOD
Lgate 1 9 1.125e-9
Ldrain 2 5 0.966e-9
Lsource 3 7 0.966e-9
RLgate 1 9 11.25
RLdrain 2 5 9.66
RLsource 3 7 9.66
Rgate 9 6 0.5
It 7 17 1
Ebreak 5 11 17 7 -550
Rbreak 17 7 RbreakMOD 1
.MODEL RbreakMOD RES (TC1=9.8e-4 TC2=-1.2e-6)
.MODEL DbodyMOD D (IS=3.9e-10  N=2.0    RS=0.209    TRS1=1.0e-4  TRS2=1.5e-7
+ CJO=3.05e-10     M=0.57      VJ=0.55  TT=3.98e-7  XTI=3        EG=1.98)
.MODEL DbreakMOD D (RS=0.1 TRS1=1e-3 TRS2=1e-6)
Rdrain 5 16 RdrainMOD 8.0
.MODEL RdrainMOD RES (TC1=7.9e-3 TC2=1.4e-5)
M_BSIM3 16 6 7 7 Bsim3 W=0.62 L=2.0e-6 NRS=1
.MODEL Bsim3 PMOS (LEVEL=7 VERSION=3.1 MOBMOD=3 CAPMOD=2 PARAMCHK=1 NQSMOD=0
+ TOX=970e-10      XJ=1.0e-6       NCH=1.3e17
+ U0=250           VSAT=5.0e5      DROUT=1.0
+ DELTA=0.1        PSCBE2=0        RSH=6.5e-3
+ VTH0=-4.00       VOFF=-0.1       NFACTOR=1.1     
+ LINT=3.45e-7     DLC=3.45e-7     CGSO=5.1e-15
+ CGSL=0           CGDO=1.2e-14    CGDL=6.65e-10
+ CJ=0             CF=0            CKAPPA=0.2
+ KT1=-1.75        KT2=0           UA1=-1.05e-9
+ NJ=10            FC=0.5)
.ends
*$
*********************** Power Discrete MOSFET Thermal Model ************************
** Product: FQB1P50
** Package: D2-PAK
**----------------------------------------------------------------------------------
.SUBCKT FQB1P50_THERMAL TH TL
CTHERM1 TH 6 2.040e-5
CTHERM2 6 5  2.180e-3
CTHERM3 5 4  8.340e-3
CTHERM4 4 3  1.620e-2
CTHERM5 3 2  2.020e-1
CTHERM6 2 TL 5.420e-1
RTHERM1 TH 6 1.300e-2
RTHERM2 6 5  2.880e-2
RTHERM3 5 4  8.680e-2
RTHERM4 4 3  4.120e-1
RTHERM5 3 2  6.580e-1
RTHERM6 2 TL 7.817e-1
.ENDS FQB1P50_THERMAL
**----------------------------------------------------------------------------------
** Creation: Mar.-24-2017   Rev.: 3.0
** ON Semiconductor
*$

